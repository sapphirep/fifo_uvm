module bindfiles;

    bind fifo fifo_assert p1 (.*);

endmodule: bindfiles