`include "fifo_base_test.sv"
`include "fifo_test1.sv"
`include "fifo_test2.sv"
`include "fifo_rand_test.sv"