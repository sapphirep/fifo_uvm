`include "fifo_base_seq.sv"
`include "fifo_seq1.sv"
`include "fifo_seq2.sv"
`include "fifo_rand_seq.sv"